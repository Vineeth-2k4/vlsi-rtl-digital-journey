module xor_gate(input A, input B, output Y);
    xor(Y, A, B);
endmodule

