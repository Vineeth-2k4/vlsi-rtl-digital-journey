module and_gate(input A, input B, output Y);
    and(Y, A, B);
endmodule


