module not_gate(input A, output Y);
    not(Y, A);
endmodule

